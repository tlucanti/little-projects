
module SN74GHC595
(

);

endmodule
